module fft016(
	f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
	f_010,f_011,f_012,f_013,f_014,f_015,
	x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
	x_010,x_011,x_012,x_013,x_014,x_015,
	W000,W001,W002,W003,W004,W005,W006,W007);
output [31:0] 
	f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
	f_010,f_011,f_012,f_013,f_014,f_015;
input [31:0] 
	x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
	x_010,x_011,x_012,x_013,x_014,x_015;
input [31:0] 
	W000,W001,W002,W003,W004,W005,W006,W007;
wire [31:0]
	x_00_000,x_00_001,x_00_002,x_00_003,x_00_004,x_00_005,x_00_006,x_00_007,x_00_008,x_00_009,
	x_00_010,x_00_011,x_00_012,x_00_013,x_00_014,x_00_015,
	x_01_000,x_01_001,x_01_002,x_01_003,x_01_004,x_01_005,x_01_006,x_01_007,x_01_008,x_01_009,
	x_01_010,x_01_011,x_01_012,x_01_013,x_01_014,x_01_015,
	x_02_000,x_02_001,x_02_002,x_02_003,x_02_004,x_02_005,x_02_006,x_02_007,x_02_008,x_02_009,
	x_02_010,x_02_011,x_02_012,x_02_013,x_02_014,x_02_015,
	x_03_000,x_03_001,x_03_002,x_03_003,x_03_004,x_03_005,x_03_006,x_03_007,x_03_008,x_03_009,
	x_03_010,x_03_011,x_03_012,x_03_013,x_03_014,x_03_015,
	x_04_000,x_04_001,x_04_002,x_04_003,x_04_004,x_04_005,x_04_006,x_04_007,x_04_008,x_04_009,
	x_04_010,x_04_011,x_04_012,x_04_013,x_04_014,x_04_015;
assign x_00_000 = x_000;
assign x_00_001 = x_001;
assign x_00_002 = x_002;
assign x_00_003 = x_003;
assign x_00_004 = x_004;
assign x_00_005 = x_005;
assign x_00_006 = x_006;
assign x_00_007 = x_007;
assign x_00_008 = x_008;
assign x_00_009 = x_009;
assign x_00_010 = x_010;
assign x_00_011 = x_011;
assign x_00_012 = x_012;
assign x_00_013 = x_013;
assign x_00_014 = x_014;
assign x_00_015 = x_015;
assign x_00_000 = x_000;
assign x_00_001 = x_001;
assign x_00_002 = x_002;
assign x_00_003 = x_003;
assign x_00_004 = x_004;
assign x_00_005 = x_005;
assign x_00_006 = x_006;
assign x_00_007 = x_007;
assign x_00_008 = x_008;
assign x_00_009 = x_009;
assign x_00_010 = x_010;
assign x_00_011 = x_011;
assign x_00_012 = x_012;
assign x_00_013 = x_013;
assign x_00_014 = x_014;
assign x_00_015 = x_015;
butt2 xx_00_000( .x0(x_00_000), .x1(x_00_008), .y0(x_01_000), .y1(x_01_008), .W(W000) );
butt2 xx_00_001( .x0(x_00_004), .x1(x_00_012), .y0(x_01_004), .y1(x_01_012), .W(W000) );
butt2 xx_00_002( .x0(x_00_002), .x1(x_00_010), .y0(x_01_002), .y1(x_01_010), .W(W000) );
butt2 xx_00_003( .x0(x_00_006), .x1(x_00_014), .y0(x_01_006), .y1(x_01_014), .W(W000) );
butt2 xx_00_004( .x0(x_00_001), .x1(x_00_009), .y0(x_01_001), .y1(x_01_009), .W(W000) );
butt2 xx_00_005( .x0(x_00_005), .x1(x_00_013), .y0(x_01_005), .y1(x_01_013), .W(W000) );
butt2 xx_00_006( .x0(x_00_003), .x1(x_00_011), .y0(x_01_003), .y1(x_01_011), .W(W000) );
butt2 xx_00_007( .x0(x_00_007), .x1(x_00_015), .y0(x_01_007), .y1(x_01_015), .W(W000) );
butt2 xx_01_000( .x0(x_01_000), .x1(x_01_004), .y0(x_02_000), .y1(x_02_004), .W(W000) );
butt2 xx_01_001( .x0(x_01_008), .x1(x_01_012), .y0(x_02_008), .y1(x_02_012), .W(W004) );
butt2 xx_01_002( .x0(x_01_002), .x1(x_01_006), .y0(x_02_002), .y1(x_02_006), .W(W000) );
butt2 xx_01_003( .x0(x_01_010), .x1(x_01_014), .y0(x_02_010), .y1(x_02_014), .W(W004) );
butt2 xx_01_004( .x0(x_01_001), .x1(x_01_005), .y0(x_02_001), .y1(x_02_005), .W(W000) );
butt2 xx_01_005( .x0(x_01_009), .x1(x_01_013), .y0(x_02_009), .y1(x_02_013), .W(W004) );
butt2 xx_01_006( .x0(x_01_003), .x1(x_01_007), .y0(x_02_003), .y1(x_02_007), .W(W000) );
butt2 xx_01_007( .x0(x_01_011), .x1(x_01_015), .y0(x_02_011), .y1(x_02_015), .W(W004) );
butt2 xx_02_000( .x0(x_02_000), .x1(x_02_002), .y0(x_03_000), .y1(x_03_002), .W(W000) );
butt2 xx_02_001( .x0(x_02_008), .x1(x_02_010), .y0(x_03_008), .y1(x_03_010), .W(W002) );
butt2 xx_02_002( .x0(x_02_004), .x1(x_02_006), .y0(x_03_004), .y1(x_03_006), .W(W004) );
butt2 xx_02_003( .x0(x_02_012), .x1(x_02_014), .y0(x_03_012), .y1(x_03_014), .W(W006) );
butt2 xx_02_004( .x0(x_02_001), .x1(x_02_003), .y0(x_03_001), .y1(x_03_003), .W(W000) );
butt2 xx_02_005( .x0(x_02_009), .x1(x_02_011), .y0(x_03_009), .y1(x_03_011), .W(W002) );
butt2 xx_02_006( .x0(x_02_005), .x1(x_02_007), .y0(x_03_005), .y1(x_03_007), .W(W004) );
butt2 xx_02_007( .x0(x_02_013), .x1(x_02_015), .y0(x_03_013), .y1(x_03_015), .W(W006) );
butt2 xx_03_000( .x0(x_03_000), .x1(x_03_001), .y0(x_04_000), .y1(x_04_001), .W(W000) );
assign f_000 = x_04_000;
assign f_008 = x_04_001;
butt2 xx_03_001( .x0(x_03_008), .x1(x_03_009), .y0(x_04_008), .y1(x_04_009), .W(W001) );
assign f_001 = x_04_008;
assign f_009 = x_04_009;
butt2 xx_03_002( .x0(x_03_004), .x1(x_03_005), .y0(x_04_004), .y1(x_04_005), .W(W002) );
assign f_002 = x_04_004;
assign f_010 = x_04_005;
butt2 xx_03_003( .x0(x_03_012), .x1(x_03_013), .y0(x_04_012), .y1(x_04_013), .W(W003) );
assign f_003 = x_04_012;
assign f_011 = x_04_013;
butt2 xx_03_004( .x0(x_03_002), .x1(x_03_003), .y0(x_04_002), .y1(x_04_003), .W(W004) );
assign f_004 = x_04_002;
assign f_012 = x_04_003;
butt2 xx_03_005( .x0(x_03_010), .x1(x_03_011), .y0(x_04_010), .y1(x_04_011), .W(W005) );
assign f_005 = x_04_010;
assign f_013 = x_04_011;
butt2 xx_03_006( .x0(x_03_006), .x1(x_03_007), .y0(x_04_006), .y1(x_04_007), .W(W006) );
assign f_006 = x_04_006;
assign f_014 = x_04_007;
butt2 xx_03_007( .x0(x_03_014), .x1(x_03_015), .y0(x_04_014), .y1(x_04_015), .W(W007) );
assign f_007 = x_04_014;
assign f_015 = x_04_015;
endmodule
////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////
module butt2(y0,y1,x0,x1,W);
  input [31:0] x0,x1,W;
  output[31:0] y0,y1;

  wire [31:0] x11;
  
  assign x11 = mulc(x1, W);
  assign y0 = addc( x0, x11 );
  assign y1 = subc( x0, x11 );
  
  function [31:0] addc;
    input [31:0] a, b;
    reg [15:0] yr, yi;
    begin
      yr = a[31:16] + b[31:16];
      yi = a[15:0] + b[15:0];
      addc = {yr, yi};
    end
  endfunction
  function [31:0] subc;
    input [31:0] a, b;
    reg [15:0] yr, yi;
    begin
      yr = a[31:16] - b[31:16];
      yi = a[15:0] - b[15:0];
      subc = {yr, yi};
    end
  endfunction
//  function [31:0] mulc;
//    input [31:0] a, b;
//    reg [15:0] yr, yi;
//    begin
//      yr = a[31:16]*b[31:16] - a[15:0]*b[15:0];
//      yi = a[15:0]*b[31:16] + a[31:16]*b[15:0];
//      mulc = {yr, yi};
//    end
//  endfunction
  function [31:0] mulc;
    input [31:0] a, b;
    reg [31:0] yr1, yr2, yi1, yi2;
    reg [15:0] ar, ai, br, bi, yyr1, yyr2, yyi1, yyi2, yr, yi;
    begin
        if( a[31] == 0 ) ar = a[31:16]; else ar = ~(a[31:16]-1);
        if( a[15] == 0 ) ai = a[15:0]; else ai = ~(a[15:0]-1);
        if( b[31] == 0 ) br = b[31:16]; else br = ~(b[31:16]-1);
        if( b[15] == 0 ) bi = b[15:0]; else bi = ~(b[15:0]-1);


        yr1 = ar * br;
        yr2 = ai * bi;

        yi1 = ar * bi;
        yi2 = ai * br;

        if( (a[31]^b[31])==0 ) yyr1 = yr1[26:11]; else yyr1 = ~yr1[26:11] + 1;
        if( (a[15]^b[15])==0 ) yyr2 = yr2[26:11]; else yyr2 = ~yr2[26:11] + 1;
        yr = yyr1 - yyr2;       

        if( (a[31]^b[15])==0 ) yyi1 = yi1[26:11]; else yyi1 = ~yi1[26:11] + 1;
        if( (a[15]^b[31])==0 ) yyi2 = yi2[26:11]; else yyi2 = ~yi2[26:11] + 1;
        yi = yyi1 + yyi2;       

      mulc = {yr, yi};
    end
  endfunction
endmodule
////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////
module top;
wire [31:0] 
	f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
	f_010,f_011,f_012,f_013,f_014,f_015;
reg [31:0] 
	x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
	x_010,x_011,x_012,x_013,x_014,x_015;
reg [31:0] 
	W000,W001,W002,W003,W004,W005,W006,W007;
fft016 f(
	f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
	f_010,f_011,f_012,f_013,f_014,f_015,
	x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
	x_010,x_011,x_012,x_013,x_014,x_015,
	W000,W001,W002,W003,W004,W005,W006,W007);
initial begin
  $dumpfile("fft.vcd");
  $dumpvars;
W000 = { 16'b 0000100000000000, 16'b 0000000000000000 };
W001 = { 16'b 0000011101100100, 16'b 1111110011110001 };
W002 = { 16'b 0000010110101000, 16'b 1111101001011000 };
W003 = { 16'b 0000001100001111, 16'b 1111100010011100 };
W004 = { 16'b 0000000000000000, 16'b 1111100000000001 };
W005 = { 16'b 1111110011110001, 16'b 1111100010011100 };
W006 = { 16'b 1111101001011000, 16'b 1111101001011000 };
W007 = { 16'b 1111100010011100, 16'b 1111110011110001 };
#100
////////
x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_001 = { 16'b 0000001111111010, 16'b 0000000000000000 };	//   0.497,  0.000
x_002 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_003 = { 16'b 0000100110011011, 16'b 0000000000000000 };	//   1.201,  0.000
x_004 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_005 = { 16'b 0000100110011011, 16'b 0000000000000000 };	//   1.201,  0.000
x_006 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_007 = { 16'b 0000001111111010, 16'b 0000000000000000 };	//   0.497,  0.000
x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_009 = { 16'b 1111110000000110, 16'b 0000000000000000 };	//  -0.497,  0.000
x_010 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_011 = { 16'b 1111011001100101, 16'b 0000000000000000 };	//  -1.201,  0.000
x_012 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_013 = { 16'b 1111011001100101, 16'b 0000000000000000 };	//  -1.201,  0.000
x_014 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_015 = { 16'b 1111110000000110, 16'b 0000000000000000 };	//  -0.497,  0.000
#100
$display( "f_000=%h", f_000);
$display( "f_001=%h", f_001);
$display( "f_002=%h", f_002);
$display( "f_003=%h", f_003);
$display( "f_004=%h", f_004);
$display( "f_005=%h", f_005);
$display( "f_006=%h", f_006);
$display( "f_007=%h", f_007);
$display( "f_008=%h", f_008);
$display( "f_009=%h", f_009);
$display( "f_010=%h", f_010);
$display( "f_011=%h", f_011);
$display( "f_012=%h", f_012);
$display( "f_013=%h", f_013);
$display( "f_014=%h", f_014);
$display( "f_015=%h", f_015);
#100
////////
x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_001 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_002 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_003 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_004 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_005 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_006 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_007 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//  -0.000,  0.000
x_009 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_010 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_011 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_012 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_013 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_014 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_015 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
#100
$display( "f_000=%h", f_000);
$display( "f_001=%h", f_001);
$display( "f_002=%h", f_002);
$display( "f_003=%h", f_003);
$display( "f_004=%h", f_004);
$display( "f_005=%h", f_005);
$display( "f_006=%h", f_006);
$display( "f_007=%h", f_007);
$display( "f_008=%h", f_008);
$display( "f_009=%h", f_009);
$display( "f_010=%h", f_010);
$display( "f_011=%h", f_011);
$display( "f_012=%h", f_012);
$display( "f_013=%h", f_013);
$display( "f_014=%h", f_014);
$display( "f_015=%h", f_015);
#100
////////
x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_001 = { 16'b 0000100110011011, 16'b 0000000000000000 };	//   1.201,  0.000
x_002 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_003 = { 16'b 1111110000000110, 16'b 0000000000000000 };	//  -0.497,  0.000
x_004 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_005 = { 16'b 1111110000000110, 16'b 0000000000000000 };	//  -0.497,  0.000
x_006 = { 16'b 0000011101011010, 16'b 0000000000000000 };	//   0.919,  0.000
x_007 = { 16'b 0000100110011011, 16'b 0000000000000000 };	//   1.201,  0.000
x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_009 = { 16'b 1111011001100101, 16'b 0000000000000000 };	//  -1.201,  0.000
x_010 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_011 = { 16'b 0000001111111010, 16'b 0000000000000000 };	//   0.497,  0.000
x_012 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_013 = { 16'b 0000001111111010, 16'b 0000000000000000 };	//   0.497,  0.000
x_014 = { 16'b 1111100010100110, 16'b 0000000000000000 };	//  -0.919,  0.000
x_015 = { 16'b 1111011001100101, 16'b 0000000000000000 };	//  -1.201,  0.000
#100
$display( "f_000=%h", f_000);
$display( "f_001=%h", f_001);
$display( "f_002=%h", f_002);
$display( "f_003=%h", f_003);
$display( "f_004=%h", f_004);
$display( "f_005=%h", f_005);
$display( "f_006=%h", f_006);
$display( "f_007=%h", f_007);
$display( "f_008=%h", f_008);
$display( "f_009=%h", f_009);
$display( "f_010=%h", f_010);
$display( "f_011=%h", f_011);
$display( "f_012=%h", f_012);
$display( "f_013=%h", f_013);
$display( "f_014=%h", f_014);
$display( "f_015=%h", f_015);
#100
////////
x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_001 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_002 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_003 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_004 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//  -0.000,  0.000
x_005 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_006 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_007 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//  -0.000,  0.000
x_009 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_010 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_011 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
x_012 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//  -0.000,  0.000
x_013 = { 16'b 0000101001100110, 16'b 0000000000000000 };	//   1.300,  0.000
x_014 = { 16'b 0000000000000000, 16'b 0000000000000000 };	//   0.000,  0.000
x_015 = { 16'b 1111010110011010, 16'b 0000000000000000 };	//  -1.300,  0.000
#100
$display( "f_000=%h", f_000);
$display( "f_001=%h", f_001);
$display( "f_002=%h", f_002);
$display( "f_003=%h", f_003);
$display( "f_004=%h", f_004);
$display( "f_005=%h", f_005);
$display( "f_006=%h", f_006);
$display( "f_007=%h", f_007);
$display( "f_008=%h", f_008);
$display( "f_009=%h", f_009);
$display( "f_010=%h", f_010);
$display( "f_011=%h", f_011);
$display( "f_012=%h", f_012);
$display( "f_013=%h", f_013);
$display( "f_014=%h", f_014);
$display( "f_015=%h", f_015);
#100
$finish;
end
endmodule
