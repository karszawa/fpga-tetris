`timescale 1ns/1ps

`define DEBUG

module tb ();

wire rst_n		;
wire sys13p5_clk	;
wire sys27_clk		;
wire sys54_clk		;
wire sys108_clk		;
wire sys100_clk	;
wire sys200_clk	;
wire sys400_clk	;
wire sys800_clk	;
wire sys120_clk	;
wire sys240_clk	;
wire sys480_clk	;
wire sys960_clk	;
wire disp40_clk	;
wire disp80_clk	;
wire disp160_clk;
wire disp320_clk;

wire sys_clk;
wire rst_sys_n;
assign sys_clk = disp40_clk;
assign rst_sys_n = rst_n;
wire disp_clk;
wire rst_disp_n;
assign disp_clk = disp40_clk;
assign rst_disp_n = rst_n;

wire        DE_OUT_HSYNC;
wire        DE_OUT_VSYNC;
wire        DE_OUT_DE;
wire [29:0] DE_OUT_RGB;

wire				clk; // 100Mhz // FPGA pin AD8
//wire				rst_n; // FPGA pin T23
wire				CLK_27MHZ_FPGA;				// FPGA pin AD13

`ifndef FOR_SIM
wire				CLK_33MHZ_FPGA; // 33Mhz // FPGA pin AB12
wire				CLK_DIFF_FPGA_P;	// E16
wire				CLK_DIFF_FPGA_N;	// E17
`else
wire				clk_40;
wire				clk_80;
wire				clk_100;
wire				clk_200;
wire				clk_120;
wire				clk_240;
wire				locked1;
wire				locked2;
`endif

	//--------------------------------------------------------------------------
	//	Chrontel 7301C Interface
	//--------------------------------------------------------------------------
wire	[11:0]		DVI_D;
wire				DVI_DE; 
wire				DVI_H; 
wire				DVI_V; 
wire				DVI_RESET_B;
wire				DVI_XCLK_P;
wire				DVI_XCLK_N; 

	//--------------------------------------------------------------------------
	//	Audio Controller in FPGA
	//--------------------------------------------------------------------------
wire				audio_bit_clk;		// FPGA pin AC13	// 12.288MHz bit clock generated by AC97
wire				audio_sdata_in;		// FPGA pin AC12	// serial data from AC97; 256bit per frame
wire				audio_sdata_out;	// FPGA pin AC11	// serial data to AC97; 256bit per frame
wire				audio_sync;			// FPGA pin AD11	// AC-Link frame sync; 12.288MHz/256 = 48kHz
wire				flash_audio_reset_b;// FPGA pin AD10	// reset of AC97; negative reset

// DIP Switches
wire	[ 8-1: 0]	DIP;

//--------------------------------------------------------------------------
//
wire				BUTTON_C; // B21
wire				BUTTON_E; // A23
wire				BUTTON_W; // C21
wire				BUTTON_S; // B22
wire				BUTTON_N; // A22

// ADC interface /* NOT USED */
wire	[ 8-1: 0]	ADN = {8{1'b0}};
wire	[ 8-1: 0]	ADP = {8{1'b1}};
wire	  			DCON= {1{1'b0}};
wire	  			DCOP= {1{1'b1}};
wire				ADC_nOE;
wire				SCLK;
wire	  			SDIO;
wire				CSB;
wire				ADCLKP;
wire				ADCLKN;

//--------------------------------------------------------------------------
// TELE_TX/RX
//--------------------------------------------------------------------------
wire				TELE_TX; // FPGA(P21 ) (HDR2_64)
wire				TELE_RX; // FPGA(AB26) (HDR1_64)
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
//	LCD Interface
//--------------------------------------------------------------------------
wire	[ 4-1: 0]	LCD_DATA	;
wire				LCD_RS		;
wire				LCD_RW		;
wire				LCD_EN  	;
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
//	I2C Bus Interface
//--------------------------------------------------------------------------
wire				I2C_SCL_DVI;
wire				I2C_SDA_DVI; 
//--------------------------------------------------------------------------
wire      			LED_C;
wire      			LED_E;
wire      			LED_W;
wire      			LED_S;
wire      			LED_N;
wire      			LED_ERR_1;
wire      			LED_ERR_0;
wire	[ 8-1: 0]	TP;


crg A0_CRG (
.rst_n			(rst_n			),//o
.sys13p5_clk	(sys13p5_clk	),//o
.sys27_clk		(sys27_clk		),//o
.sys54_clk		(sys54_clk		),//o
.sys108_clk		(sys108_clk		),//o
.sys100_clk		(sys100_clk		),//o
.sys200_clk		(sys200_clk		),//o
.sys400_clk		(sys400_clk		),//o
.sys800_clk		(sys800_clk		),//o
.sys120_clk		(sys120_clk		),//o
.sys240_clk		(sys240_clk		),//o
.sys480_clk		(sys480_clk		),//o
.sys960_clk		(sys960_clk		),//o
.disp40_clk		(disp40_clk		),//o
.disp80_clk		(disp80_clk		),//o
.disp160_clk	(disp160_clk	),//o
.disp320_clk	(disp320_clk	) //o
);


fpga_top A_FPGA_TOP (
//--------------------------------------------------------------------------
//	Clock and Reset
//--------------------------------------------------------------------------
.clk				(sys100_clk			),//i	// 100Mhz // FPGA pin AD8
.rst_n				(rst_n				),//i	// FPGA pin T23
.CLK_27MHZ_FPGA		(sys27_clk			),//i	// FPGA pin AD13
`ifndef FOR_SIM
.CLK_33MHZ_FPGA		(CLK_33MHZ_FPGA		),//i	// 33Mhz // FPGA pin AB12
.CLK_DIFF_FPGA_P	(CLK_DIFF_FPGA_P	),//i	// E16
.CLK_DIFF_FPGA_N	(CLK_DIFF_FPGA_N	),//i	// E17
`else
.clk_40				(disp40_clk			),//i
.clk_80				(disp80_clk			),//i
.clk_100			(sys100_clk			),//i
.clk_200			(sys200_clk			),//i
.clk_120			(sys120_clk			),//i
.clk_240			(sys240_clk			),//i
.locked1			(rst_n				),//i
.locked2			(rst_n				),//i
`endif
//--------------------------------------------------------------------------
//	Chrontel 7301C Interface
//--------------------------------------------------------------------------
.DVI_D				(DVI_D				),//o[11:0]
.DVI_DE				(DVI_DE				),//o
.DVI_H				(DVI_H				),//o
.DVI_V				(DVI_V				),//o
.DVI_RESET_B		(DVI_RESET_B		),//o
.DVI_XCLK_P			(DVI_XCLK_P			),//o
.DVI_XCLK_N			(DVI_XCLK_N			),//o

//--------------------------------------------------------------------------
//	Audio Controller in FPGA
//--------------------------------------------------------------------------
.audio_bit_clk		(audio_bit_clk		),//i
.audio_sdata_in		(audio_sdata_in		),//i
.audio_sdata_out	(audio_sdata_out	),//o
.audio_sync			(audio_sync			),//o
.flash_audio_reset_b(flash_audio_reset_b),//o

// DIP Switches
.DIP				({8{1'b0}}			),//i[7:0]

//--------------------------------------------------------------------------
//
.BUTTON_C			({1{1'b0}}			),//i
.BUTTON_E			({1{1'b0}}			),//i
.BUTTON_W			({1{1'b0}}			),//i
.BUTTON_S			({1{1'b0}}			),//i
.BUTTON_N			({1{1'b0}}			),//i

//	// ADC interface
//	.ADN				(ADN				),//i[7:0]
//	.ADP				(ADP				),//i[7:0]
//	.DCON				(DCON				),//i
//	.DCOP				(DCOP				),//i
//	.ADC_nOE			(ADC_nOE			),//o
//	.SCLK				(SCLK				),//o
//	.SDIO				(SDIO				),//io        
//	.CSB				(CSB				),//o
//	.ADCLKP				(ADCLKP				),//o
//	.ADCLKN				(ADCLKN				),//o

//--------------------------------------------------------------------------
// TELE_TX/RX
//--------------------------------------------------------------------------
.TELE_TX			(TELE_TX			),//o
.TELE_RX			(TELE_RX			),//i
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
//	LCD Interface
//--------------------------------------------------------------------------
.LCD_DATA			(LCD_DATA			),//io[ 4-1: 0]
.LCD_RS				(LCD_RS				),//o
.LCD_RW				(LCD_RW				),//o
.LCD_EN  			(LCD_EN  			),//o
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
//	I2C Bus Interface
//--------------------------------------------------------------------------
.I2C_SCL_DVI		(I2C_SCL_DVI		),//io
.I2C_SDA_DVI		(I2C_SDA_DVI		),//io
//--------------------------------------------------------------------------
.LED_C				(LED_C				),//o
.LED_E				(LED_E				),//o
.LED_W				(LED_W				),//o
.LED_S				(LED_S				),//o
.LED_N				(LED_N				),//o
.LED_ERR_1			(LED_ERR_1			),//o
.LED_ERR_0			(LED_ERR_0			),//o
.TP					(TP					) //o[7:0]
);

assign DE_OUT_VSYNC = A_FPGA_TOP.A_DVI_TELE_TXRX.A_DISPLAY.o_sync_va;
assign DE_OUT_HSYNC = A_FPGA_TOP.A_DVI_TELE_TXRX.A_DISPLAY.o_sync_ha;
assign DE_OUT_DE	= A_FPGA_TOP.A_DVI_TELE_TXRX.A_DISPLAY.o_sync_de;
//assign DE_OUT_RGB	={A_FPGA_TOP.A_DVI_TELE_TXRX.A_DISPLAY.o_red, 2'd0 ,
//					  A_FPGA_TOP.A_DVI_TELE_TXRX.A_DISPLAY.o_grn, 2'd0 ,
//					  A_FPGA_TOP.A_DVI_TELE_TXRX.A_DISPLAY.o_blu, 2'd0 };
assign DE_OUT_RGB	={A_FPGA_TOP.A_DVI_TELE_TXRX.Video[24-1:16], 2'd0 ,
					  A_FPGA_TOP.A_DVI_TELE_TXRX.Video[16-1: 8], 2'd0 ,
					  A_FPGA_TOP.A_DVI_TELE_TXRX.Video[ 8-1: 0], 2'd0 };

monitor_model A_DUMP (
.disp_clk		(disp80_clk		),
.rst_disp_n		(rst_n			),
.DE_OUT_VSYNC	(DE_OUT_VSYNC	),
.DE_OUT_HSYNC	(DE_OUT_HSYNC	),
.DE_OUT_DE		(DE_OUT_DE		),
.DE_OUT_RGB		(DE_OUT_RGB		)
);

endmodule

