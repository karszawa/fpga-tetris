// Audio Controlling in FPGA
//   ____________           ________
//   |          | ->->->->- |      | ->->->->- ||
//   |   FPGA   |           | AC97 |           || Audio Line In / Line Out
//   | Virtex-5 | -<-<-<-<- |      | -<-<-<-<- ||
//   ~~~~~~~~~~~~           ~~~~~~~~
//
// Access between FPGA and AC97, input: FPGA <- AC97, output: FPGA -> AC97

module audio (
	// 27Mhz Clock and Board Reset
	input				clk					,// FPGA Clock: 27Mhz
	input				rst_n				,// reset of FPGA, down:1, up:0

	// IF between AC97
	input				audio_bit_clk		,// 12.288MHz bit clock generated by AC97
	output				flash_audio_reset_b	,// reset of AC97, negative reset
	input				audio_sdata_in		,// serial data from AC97, 256bit per frame
	output				audio_sdata_out		,// serial data to AC97, 256bit per frame
	output				audio_sync			,// AC-Link frame sync, 12.288MHz/256 = 48kHz
	    
	// USER IF
	input				btn_c		,
	input				btn_n		,
	input				btn_e		,
	input				btn_s		,
	input				btn_w		,
	
	// LED OUTPUT for DEBUGGING
	output	[ 8-1: 0]	tp
);

wire	[ 8-1: 0]	tp_if;
wire	[ 8-1: 0]	tp_proc;

wire				if_Audio_sync			;
wire	[20-1: 0]	if_Audio_L				;
wire	[20-1: 0]	if_Audio_R				;
wire				proc_Audio_sync			;
wire	[20-1: 0]	proc_Audio_L			;
wire	[20-1: 0]	proc_Audio_R			;

audio_if A0_IF (
.clk					(clk					),//i
.rst_n					(rst_n					),//i
.audio_bit_clk			(audio_bit_clk			),//i
.flash_audio_reset_b	(flash_audio_reset_b	),//o
.audio_sdata_in			(audio_sdata_in			),//i
.audio_sdata_out		(audio_sdata_out		),//o
.audio_sync				(audio_sync				),//o
.btn_c					(btn_c					),//i
.btn_n					(btn_n					),//i
.btn_e					(btn_e					),//i
.btn_s					(btn_s					),//i
.btn_w					(btn_w					),//i
.oAudio_sync			(if_Audio_sync			),//o
.oAudio_L				(if_Audio_L				),//o[20-1: 0]
.oAudio_R				(if_Audio_R				),//o[20-1: 0]
.iAudio_sync			(proc_Audio_sync		),//i
.iAudio_L				(proc_Audio_L			),//i[20-1: 0]
.iAudio_R				(proc_Audio_R			),//i[20-1: 0]
.tp                     (tp_if                  ) //o[ 8-1: 0]
);

audio_proc A1_PROC (
.clk				(clk				),//i
.rst_n				(rst_n				),//i
.btn_c				(btn_c				),//i
.btn_n				(btn_n				),//i
.btn_e				(btn_e				),//i
.btn_s				(btn_s				),//i
.btn_w				(btn_w				),//i
.iAudio_sync		(if_Audio_sync		),//i
.iAudio_L			(if_Audio_L			),//i[20-1: 0]
.iAudio_R			(if_Audio_R			),//i[20-1: 0]
.oAudio_sync		(proc_Audio_sync	),//o
.oAudio_L			(proc_Audio_L		),//o[20-1: 0]
.oAudio_R			(proc_Audio_R		),//o[20-1: 0]
.tp                 (tp_proc            ) //o[ 4-1: 0]
);

assign tp = tp_if;

endmodule
