`timescale 1ns/1ns
`define USE_SYSELE

module fpga_top (
	//--------------------------------------------------------------------------
	//	Clock and Reset
	//--------------------------------------------------------------------------
	input					clk, // 100Mhz // FPGA pin AD8
	input					rst_n, // FPGA pin T23
	input					CLK_27MHZ_FPGA,				// FPGA pin AD13

`ifndef FOR_SIM
	input					CLK_33MHZ_FPGA, // 33Mhz // FPGA pin AB12
	input					CLK_DIFF_FPGA_P,	// E16
	input					CLK_DIFF_FPGA_N,	// E17
`else
	input					clk_40,
	input					clk_80,
	input					clk_100,
	input					clk_200,
	input					clk_120,
	input					clk_240,
	input					locked1,
	input					locked2,
`endif

	//--------------------------------------------------------------------------
	//	Chrontel 7301C Interface
	//--------------------------------------------------------------------------
	output	[11:0]			DVI_D,
	output					DVI_DE, 
	output					DVI_H, 
	output					DVI_V, 
	output					DVI_RESET_B,
	output					DVI_XCLK_N, DVI_XCLK_P,

	//--------------------------------------------------------------------------
	//	Audio Controller in FPGA
	//--------------------------------------------------------------------------
	input					audio_bit_clk,		// FPGA pin AC13	// 12.288MHz bit clock generated by AC97
	input					audio_sdata_in,		// FPGA pin AC12	// serial data from AC97, 256bit per frame
	output					audio_sdata_out,	// FPGA pin AC11	// serial data to AC97, 256bit per frame
	output					audio_sync,			// FPGA pin AD11	// AC-Link frame sync, 12.288MHz/256 = 48kHz
	output					flash_audio_reset_b,// FPGA pin AD10	// reset of AC97, negative reset

	// DIP Switches
	input	[7:0]			DIP,

	//--------------------------------------------------------------------------
	//
	input                   BUTTON_C, // B21
	input                   BUTTON_E, // A23
	input                   BUTTON_W, // C21
	input                   BUTTON_S, // B22
	input                   BUTTON_N, // A22

//   // ADC interface /* NOT USED */
//	input	[ 8-1: 0]		ADN,
//	input	[ 8-1: 0]		ADP,
//	input					DCON,
//	input					DCOP,
//	output					ADC_nOE,
//	output					SCLK,
//	inout					SDIO,
//	output					CSB,
//	output					ADCLKP,
//	output					ADCLKN,

	//--------------------------------------------------------------------------
	// TELE_TX/RX
	//--------------------------------------------------------------------------
	output                  TELE_TX, // FPGA(P21 ) (HDR2_64)
	input                   TELE_RX, // FPGA(AB26) (HDR1_64)
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	LCD Interface
	//--------------------------------------------------------------------------
	inout	[ 4-1: 0]		LCD_DATA	,
	output					LCD_RS		,
	output					LCD_RW		,
	output					LCD_EN  	,
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	PS/2 Interface
	//--------------------------------------------------------------------------
	inout		MOUSE_CLK		,// FPGA(L2)
	inout		MOUSE_DATA		,// FPGA(K1)
	inout		KEYBOARD_CLK	,// FPGA(J1)
	inout		KEYBOARD_DATA	,// FPGA(H2)

	//--------------------------------------------------------------------------
	//	I2C Bus Interface
	//--------------------------------------------------------------------------
	inout					I2C_SCL_DVI,
	inout					I2C_SDA_DVI, 
	//--------------------------------------------------------------------------
	output      			LED_C,
	output      			LED_E,
	output      			LED_W,
	output      			LED_S,
	output      			LED_N,
	output      			LED_ERR_1,
	output      			LED_ERR_0,
	output [7:0]			TP


);

wire	[ 8-1: 0]	TP_DVI;
wire	[ 8-1: 0]	TP_AUD;
wire	[ 8-1: 0]	TP_PS2;
wire	[ 8-1: 0]	TP_LCD;
//assign	TP = { TP_DVI[ 2-1: 0], TP_AUD[ 6-1: 0] };
//assign	TP = TP_AUD;
assign	TP = TP_LCD;

wire				mouse_valid;
wire	[12-1: 0]	mpos_x	;// current mouse position; 12 bits
wire	[12-1: 0]	mpos_y	;
wire	[ 9-1: 0]	mdif_x	;// incremental mouse position; 8 bits
wire	[ 9-1: 0]	mdif_y	;
wire				mbtn_left;
wire				mbtn_middle;
wire				mbtn_right;
wire				key_valid;
wire	[ 8-1: 0]	key_data;

`ifndef DVI_ONLY_FPGA_TOP
`ifndef FOR_SIM
wire Clock50;
wire Clock75;
wire CLKIN_IBUFG_OUT;
wire CLK0_OUT;
wire LOCKED_OUT;
crg A_CRG (
//	.CLKIN_IN(CLK_33MHZ_FPGA), 
    .CLKIN_IN(clk), 
    .RST_IN(~rst_n), 
    .CLKDV_OUT(Clock50), 
    .CLKFX_OUT(Clock75), 
    .CLKIN_IBUFG_OUT(CLKIN_IBUFG_OUT), 
    .CLK0_OUT(CLK0_OUT),
    .LOCKED_OUT(LOCKED_OUT)
);
assign clk_50 = Clock50;
assign clk_75 = Clock75;
`else //FOR_SIM
assign clk_50 = clk_80;
assign clk_75 = clk_80;
`endif //FOR_SIM
`else
`endif

DVI_TOP A_DVI_TELE_TXRX (
.clk					(clk					),//i	// 100Mhz
.rst_n					(rst_n					),//i	
`ifdef DVI_ONLY_FPGA_TOP
.CLK_33MHZ_FPGA			(CLK_33MHZ_FPGA			),//i	// 33Mhz
`else
.clk_75					(clk_75					),//i
`endif
//--------------------------------------------------------------------------
//	Chrontel 7301C Interface
//--------------------------------------------------------------------------
.DVI_D					(DVI_D					),//o[11:0]			
.DVI_DE					(DVI_DE					),//o
.DVI_H					(DVI_H					),//o
.DVI_V					(DVI_V					),//o
.DVI_RESET_B			(DVI_RESET_B			),//o
.DVI_XCLK_N				(DVI_XCLK_N				),//o
.DVI_XCLK_P				(DVI_XCLK_P				),//o
//--------------------------------------------------------------------------
//
.BUTTON_C				(BUTTON_C				),//i	// B21
.BUTTON_E				(BUTTON_E				),//i	// A23
.BUTTON_W				(BUTTON_W				),//i	// C21
.BUTTON_S				(BUTTON_S				),//i	// B22
.BUTTON_N				(BUTTON_N				),//i	// A22
.mouse_valid			(mouse_valid			),//i
.rect_pos_x				(mpos_x					),//i[12-1: 0]	
.rect_pos_y				(mpos_y					),//i[12-1: 0]	
.mouse_dif_x			(mdif_x					),//i[ 9-1: 0]	
.mouse_dif_y			(mdif_y					),//i[ 9-1: 0]	
//--------------------------------------------------------------------------
// TELE_TX/RX
//--------------------------------------------------------------------------
.TELE_TX				(TELE_TX				),//o	// P21 (HDR2_64)
.TELE_RX				(TELE_RX				),//i	// AB26(HDR1_64)
//--------------------------------------------------------------------------

`ifndef USE_SYSELE
//--------------------------------------------------------------------------
//	LCD Interface
//--------------------------------------------------------------------------
.LCD_DATA				(	{4{1'bz}}			),//io[ 4-1: 0]		
.LCD_RS					(	/* OPEN */			),//o
.LCD_RW					(	/* OPEN */			),//o
.LCD_EN  				(	/* OPEN */			),//o
//--------------------------------------------------------------------------
`endif

//--------------------------------------------------------------------------
//	I2C Bus Interface
//--------------------------------------------------------------------------
.I2C_SCL_DVI			(I2C_SCL_DVI			),//io
.I2C_SDA_DVI			(I2C_SDA_DVI			),//io
//--------------------------------------------------------------------------
.LED_C					(LED_C					),//o
.LED_E					(LED_E					),//o
.LED_W					(LED_W					),//o
.LED_S					(LED_S					),//o
.LED_N					(LED_N					),//o
.LED_ERR_1				(LED_ERR_1				),//o
.LED_ERR_0				(LED_ERR_0				),//o
.TP						(TP_DVI					) //o[7:0]
);

lcd_top A_LCD (
// Global 100MHz clock
`ifndef FOR_SIM
.CLK					(clk					),//i
.CLK50M					(clk_50					),//i
.CLK_33MHZ_FPGA			(CLK_33MHZ_FPGA			),//i
.CLK_DIFF_FPGA_P		(CLK_DIFF_FPGA_P		),//i
.CLK_DIFF_FPGA_N		(CLK_DIFF_FPGA_N		),//i
`else
.clk_40					(clk_40					),//i
.clk_100				(clk_100				),//i
.clk_200				(clk_200				),//i
.clk_120				(clk_120				),//i
.clk_240				(clk_240				),//i
.locked1				(locked1				),//i
.locked2				(locked2				),//i
`endif
// Reset signal, active low
.nRST					(rst_n					),//i
// KEYBOARD IN
.valid_i				(key_valid				),//i
.recv_data				(key_data				),//i[7:0]
// North, East, South, West and Center buttons
// Active High
.BTN_N					(BUTTON_N				),//i
.BTN_E					(BUTTON_E				),//i
.BTN_S					(BUTTON_S				),//i
.BTN_W					(BUTTON_W				),//i
.BTN_C					(BUTTON_C				),//i
// LCD driver
.LCDDATA				(LCD_DATA				),//io[3:0]
.RS						(LCD_RS					),//o
.RW						(LCD_RW					),//o
.EN						(LCD_EN  				),//o
.LED					(TP_LCD					) //o[7:0]
);


audio A_AUDIO (
.clk					(CLK_27MHZ_FPGA			),//i	// FPGA pin AD13
.rst_n					(rst_n					),//i	// FPGA pin T23		// reset of FPGA, down:1, up:0
.btn_c					(BUTTON_C				),//i
.btn_n					(BUTTON_N				),//i
.btn_e					(BUTTON_E				),//i
.btn_s					(BUTTON_S				),//i
.btn_w					(BUTTON_W				),//i
.audio_bit_clk			(audio_bit_clk			),//i	// FPGA pin AC13 (bank 4)	// 12.288MHz bit clock generated by AC97
.audio_sdata_in			(audio_sdata_in			),//i	// FPGA pin AC12 (bank 4)	// serial data from AC97, 256bit per frame
.audio_sdata_out		(audio_sdata_out		),//o	// FPGA pin AC11 (bank 4)	// serial data to AC97, 256bit per frame
.audio_sync				(audio_sync				),//o	// FPGA pin AD11 (bank 4)	// AC-Link frame sync, 12.288MHz/256 = 48kHz
.flash_audio_reset_b	(flash_audio_reset_b	),//o	// FPGA pin AD10 (bank 4)	// reset of AC97, negative reset
.tp						(TP_AUD					) //o[ 8-1: 0]
);

ps2_top A_PS2_KEY_MOUSE (
.sys50_clk				(clk_50					),//i
.rst_n					(rst_n					),//i
.MOUSE_CLK				(MOUSE_CLK				),//io
.MOUSE_DATA				(MOUSE_DATA				),//io
.KEYBOARD_CLK			(KEYBOARD_CLK			),//io
.KEYBOARD_DATA			(KEYBOARD_DATA			),//io
.mouse_valid			(mouse_valid			),//o
.mpos_x					(mpos_x					),//o[12-1: 0]	
.mpos_y					(mpos_y					),//o[12-1: 0]	
.mdif_x					(mdif_x					),//o[ 9-1: 0]	
.mdif_y					(mdif_y					),//o[ 9-1: 0]	
.mbtn_left				(mbtn_left				),//o
.mbtn_middle			(mbtn_middle			),//o
.mbtn_right				(mbtn_right				),//o
.key_valid				(key_valid				),//o
.key_data				(key_data				),//o[ 8-1: 0]	
.TP         			(TP_PS2     			) //o[ 8-1: 0]	
);

endmodule

