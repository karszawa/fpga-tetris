`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:24:48 11/30/2017 
// Design Name: 
// Module Name:    update_position 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module update_position(
    input clk,
    input i_pls_e,
    input i_pls_w,
    input board,
    input block_id,
    input block_rad,
    output blk_pos_x,
    output blk_pos_y,
    inout state
);

endmodule
